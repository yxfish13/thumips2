----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    16:02:56 11/22/2015 
-- Design Name: 
-- Module Name:    IF_inst - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity IF_inst is
    Port ( PC : in  STD_LOGIC_VECTOR (15 downto 0);
           PC_1 : out  STD_LOGIC_VECTOR (15 downto 0);
           IF_inst : out  STD_LOGIC_VECTOR (15 downto 0));
end IF_inst;

architecture Behavioral of IF_inst is

begin


end Behavioral;

